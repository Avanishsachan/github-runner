module tb;
endmodule

